----------------------------------------------------------------------------------------------------
-- PIF_RTC.vhd    pif real time clock
--
-- Initial entry: 16.06.13 sangil
--
-- Copyright (c) 2015 to 2016
--
----------------------------------------------------------------------------------------------------

----------------------------------------------------------------------------------------------------
--
----------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

----------------------------------------------------------------------------------------------------
--
----------------------------------------------------------------------------------------------------
--library work;           
--use work.defs.all;

----------------------------------------------------------------------------------------------------
--
----------------------------------------------------------------------------------------------------
--library machxo2;        
--use machxo2.components.all;

----------------------------------------------------------------------------------------------------
--
----------------------------------------------------------------------------------------------------
entity PIF_RTC is
	port 
	(	
		RST					: in std_logic;
		CLOCK				: in std_logic; -- 26.60MHz, 48.54ns
		PPS_P				: out std_logic;
		PPS_R				: out std_logic
	);
end PIF_RTC;

----------------------------------------------------------------------------------------------------
--
----------------------------------------------------------------------------------------------------
architecture rtl of PIF_RTC is

----------------------------------------------------------------------------------------------------
-- signal
----------------------------------------------------------------------------------------------------
signal pps_p_sig			: std_logic;
signal pps_r_sig			: std_logic;

----------------------------------------------------------------------------------------------------
-- constant
----------------------------------------------------------------------------------------------------
constant one_sec_period		: unsigned(23 downto 0) := "110010101111000100100000"; -- 13300000, 500ms

----------------------------------------------------------------------------------------------------
-- unsigned
----------------------------------------------------------------------------------------------------
signal one_sec_cnt			: unsigned(23 downto 0) := (others=>'0');

----------------------------------------------------------------------------------------------------
begin
----------------------------------------------------------------------------------------------------
PPS_P <= pps_p_sig;
PPS_R <= pps_r_sig;

process(RST, CLOCK)
begin
	if (RST = '0') then
		one_sec_cnt <= (others => '0');
		pps_p_sig <= '0';
		pps_r_sig <= '0';
	elsif rising_edge(CLOCK) then
		one_sec_cnt <= one_sec_cnt + 1;
		if (one_sec_cnt = one_sec_period) then -- 500 ms
			pps_p_sig <= not pps_p_sig;
			pps_r_sig <= not pps_r_sig;
			one_sec_cnt <= (others => '0');
		end if;
	end if;
end process;

----------------------------------------------------------------------------------------------------
end rtl;
----------------------------------------------------------------------------------------------------